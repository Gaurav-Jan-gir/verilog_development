module andGate (A, B, C);
    input A, B;
    output C;

    assign C = A & B; // AND operation
endmodule
// Testbench for the AND gate