module xorGate(A,B,C);
    input A, B;
    output C;

    assign C = A ^ B; // XOR operation
endmodule