module orGate (A, B, Y);
    input A, B;
    output Y;
    
    assign Y = A | B; // OR operation
endmodule
